package ca12_dat_103 is

constant ca12_type103:integer:=1;
constant ca12_inve103:integer:=2;
signal ca12_ord103:real_vector(1 to 3):=(6.0, 2.0, 0.0);
signal ca12_fak103:real_vector(1 to 4):=(0.340259232109, 8.27974055976, 0.00000000000, 462.927518575);
constant ca12_anz103:integer:=       21;
signal ca12_data103:real_vector(1 to 21):=
(
  0.753283687900    ,
  0.274473414578    ,
 -0.461863149061E-01,
  0.138701246697E-01,
 -0.577173008909E-02,
  0.872396318797E-02,
 -0.551446912259E-02,
  0.497764560409E-02,
  0.375266194850E-02,
 -0.237433276804E-02,
  0.793317695316E-03,
 -0.345447049565E-03,
  0.181030057463E-02,
 -0.135055776377E-02,
 -0.240462928166E-03,
  0.174907882002E-03,
 -0.150577377133E-03,
 -0.372662233549E-04,
  0.721515427319E-04,
  0.276041714666E-03,
 -0.246811712009E-03
);
end;
