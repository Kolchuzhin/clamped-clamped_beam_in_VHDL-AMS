package s_dat_103 is

constant s_type103:integer:=1;
constant s_inve103:integer:=1;
signal s_ord103:real_vector(1 to 3):=( 6.0    , 2.0    , 0.0    );
signal s_fak103:real_vector(1 to 4):=(  0.340259232109    ,   8.27974055976    ,   0.00000000000    ,   2338.04387300    );
constant s_anz103:integer:=      21;
signal s_data103:real_vector(1 to       21):=
(
  0.246103007688E-01,
 -0.592194289171E-14,
  0.588163120255    ,
  0.206195084844E-13,
  0.310785053702    ,
 -0.150090189401E-13,
  0.218511103401E-03,
  0.561671007347E-16,
 -0.607923437658E-03,
 -0.974081033856E-15,
 -0.397309376326E-01,
  0.253061854361E-14,
 -0.177980113126E-04,
 -0.162208591397E-14,
  0.253678100458E-01,
  0.691613737529E-14,
  0.104640619917E-01,
 -0.245661412821E-13,
  0.344132820990E-04,
  0.180081497945E-13,
  0.700669792426E-07
);
end;
