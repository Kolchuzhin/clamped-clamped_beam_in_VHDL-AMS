package initial is

constant mm_1:real:= 0.185207030268E-11;
constant dm_1:real:= 0.00000000000 ;
constant mm_2:real:= 0.194379055271E-11;
constant dm_2:real:= 0.00000000000 ;
constant fi1_1:real:= 0.995464482369 ;
constant fi1_2:real:= -0.929504617585 ;
constant fi2_1:real:= 0.553419215537 ;
constant fi2_2:real:= 0.888589814646 ;
constant el1_1:real:= -24.1171438098 ;
constant el1_2:real:= -10.6523772382 ;
constant el2_1:real:= 52.6096410185 ;
constant el2_2:real:= 23.3814480531 ;

end;
